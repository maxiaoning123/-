module Bluetooth_dataa(
    input                     clk,
    input                     rst_n,
    input   [31:0]            duty_cycle/* synthesis PAP_MARK_DEBUG="1"*/,  // ռ�ձȣ�0-100��
    input   [19:0]            ad_fred/* synthesis PAP_MARK_DEBUG="1"*/,     // Ƶ�ʣ�0-1048575��
    input   [7:0]             ad_max/* synthesis PAP_MARK_DEBUG="1"*/,      // ADC��������128-255��
	 
    input                     uart_tx_done, // UART��������ź�
    input   [7:0]             uart_rx_data, // UART��������
    input                     uart_rx_done, // UART��������ź�
    
    output  reg               uart_tx_en/* synthesis PAP_MARK_DEBUG="1"*/,   // UART����ʹ��
    output  reg     [7:0]     uart_tx_data/* synthesis PAP_MARK_DEBUG="1"*/   // UART��������
    

);
	 
// ״̬����
parameter IDLE              = 4'd0;  // ����̬
parameter DATA_CHANGE       = 4'd1;  // ���ݷֽ�����Чλ�滻̬
parameter WAIT_1s           = 4'd2;  // �ȴ�1s
parameter SEND              = 4'd3;  // UART����̬
parameter OVER              = 4'd4;  // �������̬

// �ȴ�1s�������ֵ
parameter count_max         = 32'd50_000_000;
reg  [7:0]   max_tx_count/* synthesis PAP_MARK_DEBUG="1"*/;  // �����ݷ����ֽ�����duty:12, fred:16, mv:13��

reg [15:0]        ad_mv_output; // 16λģ���ֵ���

// ״̬��������Ĵ���
reg  [3:0]    state/* synthesis PAP_MARK_DEBUG="1"*/;        // ��ǰ״̬
reg  [31:0]   count;        // WAIT_1s����
reg  [5:0]    tx_count/* synthesis PAP_MARK_DEBUG="1"*/;     // �����ֽڼ���
reg  [1:0]    tx_en_count;  // ����ʹ�ܼ���
reg           uart_tx_en_temp; // ����ʹ����ʱ�ź�
reg  [1:0]    change_count/* synthesis PAP_MARK_DEBUG="1"*/; // �����л�������0:duty,1:fred,2:mv��

// -------------------------- 1. ���ݷֽ�����Чλ�滻�����߼� --------------------------
// 1.1 ԭʼASCII�ֽ�Ĵ�������ʱ�洢δ�����ASCII�룩
reg [7:0] duty_ascii_raw [2:0];  // ռ�ձ�ԭʼASCII
reg [7:0] fred_ascii_raw [6:0];  // Ƶ��ԭʼASCII
reg [7:0] mv_ascii_raw [4:0];    // ģ���ֵԭʼASCII��[4]��λ,[3]ǧλ,[2]��λ,[1]ʮλ,[0]��λ (5λ, max 49784)

// 1.2 ���շ���ASCII�Ĵ�������Чλ���滻Ϊ�ո�
reg [7:0] duty_ascii_final [2:0]; // ռ�ձ�����ASCII
reg [7:0] fred_ascii_final [6:0]; // Ƶ������ASCII
reg [7:0] mv_ascii_final [4:0];   // ģ���ֵ����ASCII

// 1.3 ��ʱ���ݼĴ������洢�޷�������ݣ�
reg [31:0] temp_duty;  // �޷���ռ�ձȣ�0-100��
reg [19:0] temp_fred;  // Ƶ�ʣ�0-1048575��
reg [15:0] ad_mv;      // 16λ�޷���ģ���ֵ��0-49784��
reg [8:0]  ad_max_minus_128; // 9λ�޷���������� 255-128 = 127

// -------------------------- 2. ����1��ԭʼ���ݷֽ⣨ת��ΪASCII�� --------------------------
// 2.1 ռ�ձȷֽ⣨ԭ�߼����䣩
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        temp_duty <= 32'd0;
        duty_ascii_raw[0] <= 8'h30;
        duty_ascii_raw[1] <= 8'h30;
        duty_ascii_raw[2] <= 8'h30;
    end
    else begin
        // ռ�ձ��޷�������0-100���߽紦��
        temp_duty <= (duty_cycle > 1000) ? 32'd999 : (duty_cycle < 0 ? 32'd0 : duty_cycle);
        // ת��ΪASCII��0��8'h30��9��8'h39��
        duty_ascii_raw[0] <= (temp_duty % 10) + 8'h30;        // ��λ
        duty_ascii_raw[1] <= ((temp_duty % 100) / 10) + 8'h30;// ʮλ
        duty_ascii_raw[2] <= (temp_duty / 100) + 8'h30;       // ��λ
    end
end

// 2.2 Ƶ�ʷֽ⣨ԭ�߼����䣩
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        temp_fred <= 20'd0;
        fred_ascii_raw[0] <= 8'h30;
        fred_ascii_raw[1] <= 8'h30;
        fred_ascii_raw[2] <= 8'h30;
        fred_ascii_raw[3] <= 8'h30;
        fred_ascii_raw[4] <= 8'h30;
        fred_ascii_raw[5] <= 8'h30;
        fred_ascii_raw[6] <= 8'h30;
    end
    else begin
        temp_fred <= ad_fred;
        // ת��ΪASCII
        fred_ascii_raw[0] <= (temp_fred / 1000000) + 8'h30;        // ����λ
        fred_ascii_raw[1] <= ((temp_fred % 1000000) / 100000) + 8'h30;// ʮ��λ
        fred_ascii_raw[2] <= ((temp_fred % 100000) / 10000) + 8'h30;  // ��λ
        fred_ascii_raw[3] <= ((temp_fred % 10000) / 1000) + 8'h30;    // ǧλ
        fred_ascii_raw[4] <= ((temp_fred % 1000) / 100) + 8'h30;     // ��λ
        fred_ascii_raw[5] <= ((temp_fred % 100) / 10) + 8'h30;       // ʮλ
        fred_ascii_raw[6] <= (temp_fred % 10) + 8'h30;               // ��λ
    end
end

// 2.3 ģ���ֵ ad_mv ����ͷֽ� (�滻ԭad_max�ֽ��߼�)
always @(posedge clk or negedge rst_n) begin
    
    
    if (!rst_n) begin
        ad_mv <= 16'd0;
        mv_ascii_raw[0] <= 8'h30;
        mv_ascii_raw[1] <= 8'h30;
        mv_ascii_raw[2] <= 8'h30;
        mv_ascii_raw[3] <= 8'h30;
        mv_ascii_raw[4] <= 8'h30;
        ad_mv_output <= 16'd0;
    end
    else begin
        // ���� ad_mv = (ad_max - 128) * 392
        // ���� ad_max ��Χ [128, 255]�� ad_max - 128 ��Χ [0, 127]
        ad_max_minus_128 <= ad_max - 8'd128; // ȷ�� ad_max ��С�� 128
        
        // 16'd392 * 9'd127 = 49784 < 65536�� 16λ�޷������㹻
        ad_mv <= ad_max_minus_128 * 16'd392; 
        ad_mv_output <= ad_mv; // �������
        
        // ת��ΪASCII (5λ���֣����49784)
        mv_ascii_raw[0] <= (ad_mv % 10) + 8'h30;          // ��λ
        mv_ascii_raw[1] <= ((ad_mv / 10) % 10) + 8'h30;   // ʮλ
        mv_ascii_raw[2] <= ((ad_mv / 100) % 10) + 8'h30;  // ��λ
        mv_ascii_raw[3] <= ((ad_mv / 1000) % 10) + 8'h30; // ǧλ
        mv_ascii_raw[4] <= (ad_mv / 10000) + 8'h30;       // ��λ
    end
end


// -------------------------- 3. ����2����Чλ�滻 --------------------------
// 3.1 ռ�ձ���Чλ�滻��ԭ�߼����䣩
always @(*) begin
    if (!rst_n) begin
        duty_ascii_final[0] = 8'h30;
        duty_ascii_final[1] = 8'h30;
        duty_ascii_final[2] = 8'h30;
    end
    else begin
        // ... (ԭռ�ձ���Чλ�滻�߼�) ...
        duty_ascii_final[0] = duty_ascii_raw[0];
        
        if (temp_duty < 10 && duty_ascii_raw[2] == 8'h30) 
            duty_ascii_final[1] = 8'h20; // �ո�
        else 
            duty_ascii_final[1] = duty_ascii_raw[1];
        
        if (temp_duty < 100) 
            duty_ascii_final[2] = 8'h20; // �ո�
        else 
            duty_ascii_final[2] = duty_ascii_raw[2];
    end
end

// 3.2 Ƶ����Чλ�滻��ԭ�߼����䣩
always @(*) begin
    if (!rst_n) begin
        // ... (��λ״̬) ...
        fred_ascii_final[0] = 8'h30;
        fred_ascii_final[1] = 8'h30;
        fred_ascii_final[2] = 8'h30;
        fred_ascii_final[3] = 8'h30;
        fred_ascii_final[4] = 8'h30;
        fred_ascii_final[5] = 8'h30;
        fred_ascii_final[6] = 8'h30;
    end
    else begin
        // ... (ԭƵ����Чλ�滻�߼�) ...
        fred_ascii_final[6] = fred_ascii_raw[6];
        
        if (temp_fred < 10 && (fred_ascii_raw[0] == 8'h30) && (fred_ascii_raw[1] == 8'h30) 
            && (fred_ascii_raw[2] == 8'h30) && (fred_ascii_raw[3] == 8'h30) && (fred_ascii_raw[4] == 8'h30))
            fred_ascii_final[5] = 8'h20;
        else
            fred_ascii_final[5] = fred_ascii_raw[5];
        
        if (temp_fred < 100 && (fred_ascii_raw[0] == 8'h30) && (fred_ascii_raw[1] == 8'h30) 
            && (fred_ascii_raw[2] == 8'h30) && (fred_ascii_raw[3] == 8'h30))
            fred_ascii_final[4] = 8'h20;
        else
            fred_ascii_final[4] = fred_ascii_raw[4];
        
        if (temp_fred < 1000 && (fred_ascii_raw[0] == 8'h30) && (fred_ascii_raw[1] == 8'h30) && (fred_ascii_raw[2] == 8'h30))
            fred_ascii_final[3] = 8'h20;
        else
            fred_ascii_final[3] = fred_ascii_raw[3];
        
        if (temp_fred < 10000 && (fred_ascii_raw[0] == 8'h30) && (fred_ascii_raw[1] == 8'h30))
            fred_ascii_final[2] = 8'h20;
        else
            fred_ascii_final[2] = fred_ascii_raw[2];
        
        if (temp_fred < 100000 && (fred_ascii_raw[0] == 8'h30))
            fred_ascii_final[1] = 8'h20;
        else
            fred_ascii_final[1] = fred_ascii_raw[1];
        
        if (temp_fred < 1000000)
            fred_ascii_final[0] = 8'h20;
        else
            fred_ascii_final[0] = fred_ascii_raw[0];
    end
end

// 3.3 ģ���ֵ ad_mv ��Чλ�滻���滻ԭad_max�߼���
always @(*) begin
    if (!rst_n) begin
        mv_ascii_final[0] = 8'h30;
        mv_ascii_final[1] = 8'h30;
        mv_ascii_final[2] = 8'h30;
        mv_ascii_final[3] = 8'h30;
        mv_ascii_final[4] = 8'h30;
    end
    else begin
        // ��λ��ʼ����Ч
        mv_ascii_final[0] = mv_ascii_raw[0];
        
        // ʮλ������"���ݣ�10"ʱ��Ч
        if (ad_mv < 10) 
            mv_ascii_final[1] = 8'h20; // �ո�
        else 
            mv_ascii_final[1] = mv_ascii_raw[1];
        
        // ��λ������"���ݣ�100"ʱ��Ч
        if (ad_mv < 100) 
            mv_ascii_final[2] = 8'h20; // �ո�
        else 
            mv_ascii_final[2] = mv_ascii_raw[2];
        
        // ǧλ������"���ݣ�1000"ʱ��Ч
        if (ad_mv < 1000) 
            mv_ascii_final[3] = 8'h20; // �ո�
        else 
            mv_ascii_final[3] = mv_ascii_raw[3];
        
        // ��λ������"���ݣ�10000"ʱ��Ч
        if (ad_mv < 10000) 
            mv_ascii_final[4] = 8'h20; // �ո�
        else 
            mv_ascii_final[4] = mv_ascii_raw[4];
    end
end


// -------------------------- 4. ����3��UART��������ѡ�� --------------------------
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        uart_tx_data <= 8'd0;
    end
    // ����ռ�ձȣ�change_count=0��
    else if (change_count == 2'd0 && state == SEND) begin
        case(tx_count)
            6'd0: uart_tx_data <= 8'h64; // "d"
            6'd1: uart_tx_data <= 8'h75; // "u"
            6'd2: uart_tx_data <= 8'h74; // "t"
            6'd3: uart_tx_data <= 8'h79; // "y"
            6'd4: uart_tx_data <= 8'h3A; // ":"
            6'd5: uart_tx_data <= duty_ascii_final[2];
            6'd6: uart_tx_data <= duty_ascii_final[1];
            6'd7: uart_tx_data <= 8'h2E; // "."
            6'd8: uart_tx_data <= duty_ascii_final[0];
            6'd9: uart_tx_data <= 8'h25; // "%"
            6'd10: uart_tx_data <= 8'h0D; // "\r"
            6'd11:uart_tx_data <= 8'h0A; // "\n"
            default: uart_tx_data <= 8'd0;
        endcase
    end
    // ����Ƶ�ʣ�change_count=1��
    else if (change_count == 2'd1 && state == SEND) begin
        case(tx_count)
            6'd0: uart_tx_data <= 8'h66; // "f"
            6'd1: uart_tx_data <= 8'h72; // "r"
            6'd2: uart_tx_data <= 8'h65; // "e"
            6'd3: uart_tx_data <= 8'h71; // "q"
            6'd4: uart_tx_data <= 8'h3A; // ":"
            6'd5: uart_tx_data <= fred_ascii_final[0];
            6'd6: uart_tx_data <= fred_ascii_final[1];
            6'd7: uart_tx_data <= fred_ascii_final[2];
            6'd8: uart_tx_data <= fred_ascii_final[3];
            6'd9: uart_tx_data <= fred_ascii_final[4];
            6'd10:uart_tx_data <= fred_ascii_final[5];
            6'd11:uart_tx_data <= fred_ascii_final[6];
            6'd12:uart_tx_data <= 8'h48; // "H"
            6'd13:uart_tx_data <= 8'h7A; // "z"
            6'd14:uart_tx_data <= 8'h0D; // "\r"
            6'd15:uart_tx_data <= 8'h0A; // "\n"
            default: uart_tx_data <= 8'd0;
        endcase
    end
    // ����ģ���ֵ ad_mv��change_count=2��(�µ��߼�)
    else if (change_count == 2'd2 && state == SEND) begin
        case(tx_count)
            6'd0: uart_tx_data <= 8'h61; // "a"
            6'd1: uart_tx_data <= 8'h64; // "d"
            6'd2: uart_tx_data <= 8'h6D; // "m"
            6'd3: uart_tx_data <= 8'h61; // "a"
            6'd4: uart_tx_data <= 8'h78; // "x"
            6'd5: uart_tx_data <= 8'h3A; // ":"
            6'd6: uart_tx_data <= mv_ascii_final[4]; // ��λ����Ч/�ո�
            6'd7: uart_tx_data <= mv_ascii_final[3]; // ǧλ����Ч/�ո�
            6'd8: uart_tx_data <= mv_ascii_final[2]; // ��λ����Ч/�ո�
            6'd9: uart_tx_data <= mv_ascii_final[1]; // ʮλ����Ч/�ո�
            6'd10:uart_tx_data <= 8'h20; // ��λ����Ч��
            6'd11:uart_tx_data <= 8'h6D; // "m"
            6'd12:uart_tx_data <= 8'h76; // "v"
            6'd13:uart_tx_data <= 8'h0D; // "\r"
            6'd14:uart_tx_data <= 8'h0A; // "\n"
            default: uart_tx_data <= 8'd0;
        endcase
    end
end


// -------------------------- 5. ����ʹ�ܿ��ƣ�ԭ�߼����䣩 --------------------------
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        tx_en_count <= 2'b0;
    end
    else if (state == SEND && tx_en_count < 2'd1 && tx_count == 8'd0) begin
        tx_en_count <= tx_en_count + 1'd1;
    end
    else if (state == SEND && tx_en_count == 2'd1 && tx_count == 8'd0) begin
        tx_en_count <= 2'd3;
    end
    else if (state == OVER) begin
        tx_en_count <= 2'd0;
    end
end

// -------------------------- 6. �����ֽڼ�����ԭ�߼����䣩 --------------------------
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        tx_count <= 8'd0;
    end
    else if (state == SEND && uart_tx_done == 1'd1) begin
        tx_count <= tx_count + 1'b1;
    end
    else if (state != SEND) begin
        tx_count <= 8'd0;
    end
end

// -------------------------- 7. UART����ʹ�������ԭ�߼����䣩 --------------------------
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        uart_tx_en_temp <= 1'b0;
    end
    else if (state == SEND && tx_en_count == 2'd1) begin
        uart_tx_en_temp <= 1'b1;
    end
    else if (state == SEND && tx_count < (max_tx_count - 1) && uart_tx_done == 1'd1) begin
        uart_tx_en_temp <= 1'b1;
    end
    else begin
        uart_tx_en_temp <= 1'b0;
    end
end

always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        uart_tx_en <= 1'b0;
    end
    else begin
        uart_tx_en <= uart_tx_en_temp;
    end
end

// -------------------------- 8. WAIT_1s������ԭ�߼����䣩 --------------------------
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        count <= 32'd0;
    end
    else if (state == WAIT_1s && count < count_max) begin
        count <= count + 32'd1;
    end
    else if (state == WAIT_1s && count == count_max) begin
        count <= 32'd0;
    end
end

// -------------------------- 9. ״̬����ת��ԭ�߼����䣩 --------------------------
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        state <= IDLE;
        change_count <= 2'd0;
    end
    else begin
        case(state)
            IDLE: begin
                state <= DATA_CHANGE;
            end
            DATA_CHANGE: begin
                state <= WAIT_1s;
            end
            WAIT_1s: begin
                if (count == count_max) begin
                    state <= SEND;
                end
            end
            SEND: begin
                if (tx_count == max_tx_count) begin
                    state <= OVER;
                end
            end
            OVER: begin
                state <= IDLE;
                // �л���һ�����ݣ�0:duty��1:fred��2:mv��0:dutyѭ����
                if (change_count == 2'd0) begin
                    change_count <= 2'd1;
                end
                else if (change_count == 2'd1) begin
                    change_count <= 2'd2;
                end
                else begin // change_count == 2'd2
                    change_count <= 2'd0;
                end
            end
            default: state <= IDLE;
        endcase
    end
end

// -------------------------- 10. �����ݷ����ֽ������ã����޸ģ� --------------------------
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        max_tx_count <= 8'd12;
    end
    else if (change_count == 2'd2 ) begin
        max_tx_count <= 8'd15; // ģ���ֵ ad_mv��15�ֽ�
    end
    else if (change_count == 2'd0 ) begin
        max_tx_count <= 8'd12; // ռ�ձȣ�12�ֽ�
    end
    else begin
        max_tx_count <= 8'd16; // Ƶ�ʣ�16�ֽ�
    end
end

endmodule