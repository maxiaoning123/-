module uart_data_check(
    input         clk,
    input         rst_n,
    input         uart_rx_done,   // UART ���������������Ч�ı�־��ͨ���ǵ��������壩
    input  [7:0]  uart_rx_data,   // ���յ��� 8 λ����
    
    output        Goal_inc,       // Ŀ��Ƶ���������� (��Ӧ���� '2B')
    output        Goal_dec        // Ŀ��Ƶ�ʼ�С���� (��Ӧ���� '2D')
   );

// ------------------------------------------
// I. ��������
// ------------------------------------------
// ASCII �� '2B' �� '2D'
// ע�⣺�������UART���͵���ASCII�ַ� '2' �� 'B'�������ǲ���һ���ֽ� '2B'H��
// �������� '2B' �� '2D' ��һ�����ֽڵ�ʮ������ֵ��
localparam DATA_INC = 8'h2B; // ��Ӧ Goal_inc �������ֽ�
localparam DATA_DEC = 8'h2D; // ��Ӧ Goal_dec �������ֽ�

reg r_Goal_inc;
reg r_Goal_dec;

always @(posedge clk or negedge rst_n) begin
    if (rst_n == 1'b0) begin
        r_Goal_inc <= 1'b0;
        r_Goal_dec <= 1'b0;
    end else begin
        // Goal_inc ����
        if (uart_rx_done & (uart_rx_data == DATA_INC)) begin
            r_Goal_inc <= 1'b1; // �����ݽ�����ɵ������ø�
        end else begin
            r_Goal_inc <= 1'b0; // �����õ�
        end
        
        // Goal_dec ����
        if (uart_rx_done & (uart_rx_data == DATA_DEC)) begin
            r_Goal_dec <= 1'b1; // �����ݽ�����ɵ������ø�
        end else begin
            r_Goal_dec <= 1'b0; // �����õ�
        end
    end
end

assign Goal_inc = r_Goal_inc;
assign Goal_dec = r_Goal_dec;


endmodule