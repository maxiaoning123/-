module Bluetooth_send(
    input                     sys_clk  ,  
    input                     rst_n,
       
    input            		  uart_rxd ,   
    output           		  uart_txd ,
    output                    Goal_inc ,      
    output                    Goal_dec ,      
    
    input   [31:0]            duty_cycle,
    input   [19:0]            ad_fred,
    input   [7 :0]            ad_max
    );
//uart
wire            uart_tx_en; 
wire            uart_rx_done; 
wire            uart_tx_done; 
wire  [7:0]     uart_tx_data; 
wire  [7:0]     uart_rx_data; 


uart_top uart_top_inst (
    .sys_clk      (sys_clk),    // ϵͳʱ�ӣ����� UART �ڲ�����������
    .sys_rst_n    (rst_n),        // ϵͳ��λ���͵�ƽ��Ч����ģ�鶨��һ�£�
    
    .uart_rxd     (uart_rxd), // �����ⲿ UART ��������
    .uart_txd     (uart_txd), // �����ⲿ UART ��������
    
    .uart_tx_en   (uart_tx_en),   
    .uart_rx_done (uart_rx_done), 
    .uart_tx_done (uart_tx_done), 
    
    .uart_tx_data (uart_tx_data), 
    .uart_rx_data (uart_rx_data)  
);

Bluetooth_dataa bluetooth_dataa_inst (
    .clk          (sys_clk),  // ϵͳʱ�ӣ�����UART����������
    .rst_n        (rst_n),      // ϵͳ��λ������Ч��
    
    // �����͵�ԭʼ����
    .duty_cycle   (duty_cycle),     // ռ�ձȣ�31λ��ʵ����Ч0-100��
    .ad_fred      (ad_fred),        // Ƶ�ʣ�19λ��ʵ����Ч0-9999999��
    .ad_max       (ad_max),         // ��ֵ��7λ��ʵ����Ч0-999��
    
    .uart_tx_done (uart_tx_done),   // UART������ɱ�־
    .uart_rx_data (uart_rx_data),   // UART���յ�������
    .uart_rx_done (uart_rx_done),   // UART������ɱ�־
    
    .uart_tx_en   (uart_tx_en),     // ����ʹ���ź�
    .uart_tx_data (uart_tx_data)    // �����͵��ֽ�����
);

// ----------------------------------------------------
// uart_data_check ������������
// ----------------------------------------------------
uart_data_check u_uart_decoder (
    .clk          ( sys_clk        ), // ���룺ϵͳʱ��
    .rst_n        ( rst_n      ), // ���룺��λ�ź� (����Ч)
    .uart_rx_done ( uart_rx_done     ), // ���룺UART�������/������Ч�ź�
    .uart_rx_data ( uart_rx_data ), // ���룺UART���յ���8λ���� [7:0]
    
    .Goal_inc     ( Goal_inc ), // �����Ƶ����������
    .Goal_dec     ( Goal_dec )  // �����Ƶ�ʼ�С����
);




endmodule
