`timescale 1ns/1ps 
module tb_top();

// �����źŶ���
reg         clk_27M;  // 50MHzʱ��
reg         rst_n;    // ��λ�źţ��͵�ƽ��Ч��

// ʵ��������ģ��
top u_top(
    .clk_27M  (clk_27M),
    .rst_n    (rst_n)
);


// ����50MHzʱ�ӣ�����20ns��
initial begin
    clk_27M = 1'b0;
    forever #18.52 clk_27M = ~clk_27M;  // ÿ10ns��תһ�Σ�Ƶ��50MHz
end

// ���ɸ�λ�źţ���ʼ��λ��һ��ʱ����ͷţ�
initial begin
    rst_n = 1'b0;          // ��ʼ��λ��Ч
    #100;                  // ���ָ�λ100ns
    rst_n = 1'b1;          // �ͷŸ�λ
    #100000;               // �����㹻��ʱ�䣨100us����ȷ�������ȶ�

end

GTP_GRS GRS_INST(.GRS_N (1'b1));

endmodule