/*
 * ģ��: bluetooth_data
 * ����:
 * 1. ͨ��FIFO��������ADʱ�����FFT���ݡ�
 * 2. ʹ��ϵͳʱ�� (clk) ���FSM������״̬������ȡFIFO��
 * 3. �ڷ���2048��FFT���ݵ�֮ǰ�����ȷ��������ֽڵ�֡ͷ (8'h05, 8'h64)��
 * 4. ͨ�� uart_tx_en �� uart_tx_data ����UARTģ����з��͡�
 * 5. ��2048�����ݷ�����ɺ����� uart_fft_over �źš�
 */
module bluetooth_data(
    input        clk,            // ϵͳʱ�� (����FSM��FIFO��)
    input        ad_clk,         // ADCʱ�� (����FIFOд)
    input        rst_n,          // �첽��λ (����Ч)
    input[7:0]   fft_data,       // FFT��������
    input        fft_data_vaild, // FFT������Ч�ź�
    input        uart_tx_done,   // UARTģ�鷢���������
    
    output reg   uart_tx_en,     // UART����ʹ�� (����)
    output [7:0] uart_tx_data,   // ���͸�UART������ (֡ͷ��FFT����)
    output reg   uart_fft_over     // һ֡(2048��)���ݷ�����ɱ�־
   );
   
// ----------------------------------------------------------------
// FIFO ʵ���� (�첽FIFO)
// ----------------------------------------------------------------

// FIFO �ڲ��ź�
wire        wr_full;
wire        almost_full;

reg         rd_en;          // FIFO ��ʹ�� (��FSM����)
wire[7:0]   rd_data;        // ��FIFO����������
wire        rd_empty;       // FIFO �ձ�־
wire        almost_empty;

// ʵ����FIFO (������������Ϊ 'fifo' ��IP�˻�ģ��)
fifo u_fifo (
  .wr_clk(ad_clk),                    // дʱ�� (ADCʱ����)
  .wr_rst(~rst_n),                    // д��λ (����Ч)
  .wr_en(fft_data_vaild),             // дʹ��
  .wr_data(fft_data),                 // д������
  .wr_full(wr_full),                  // output
  .almost_full(almost_full),          // output
  
  .rd_clk(clk),                       // ��ʱ�� (ϵͳʱ����)
  .rd_rst(~rst_n),                    // ����λ (����Ч)
  .rd_en(rd_en),                      // ��ʹ��
  .rd_data(rd_data),                  // ��������
  .rd_empty(rd_empty),                // output
  .almost_empty(almost_empty)         // output
);

// ----------------------------------------------------------------
// ���ڷ���FSM (����״̬��)
// ----------------------------------------------------------------

// FSM ״̬����
localparam S_IDLE         = 4'd0; // ����״̬
localparam S_SEND_HEADER1 = 4'd1; // ����֡ͷ1 (0x05)
localparam S_WAIT_HEADER1 = 4'd2; // �ȴ�֡ͷ1�������
localparam S_SEND_HEADER2 = 4'd3; // ����֡ͷ2 (0x64)
localparam S_WAIT_HEADER2 = 4'd4; // �ȴ�֡ͷ2�������
localparam S_READ_FIFO    = 4'd5; // ��FIFO��ȡ����
localparam S_SEND_UART    = 4'd6; // ����FIFO���ݵ�UART
localparam S_WAIT_UART    = 4'd7; // �ȴ�UART���ݷ������
localparam S_FINISH       = 4'd8; // 2048��ȫ���������

// FSM ״̬�Ĵ���
reg [3:0] state_reg; 
// FFT���ݷ��ͼ����� (0 �� 2047)
reg [10:0] count_reg;

// ���ڱ���֡ͷ���ݵı���
reg [7:0] header_data_reg;

// ----------------------------------------------------------------
// ����·�� MUX (����ѡ����)
// ----------------------------------------------------------------
// ����FSM״̬���� uart_tx_data �����
// ״̬ <= S_WAIT_HEADER2 (4) ʱ, ���֡ͷ
// ״̬ >  S_WAIT_HEADER2 (4) ʱ, ���FIFO����
assign uart_tx_data = (state_reg > S_WAIT_HEADER2) ? rd_data : header_data_reg;


// ----------------------------------------------------------------
// FSM �����߼� (ʱ���߼�)
// ----------------------------------------------------------------
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        // �첽��λ
        state_reg       <= S_IDLE;
        count_reg       <= 11'd0;
        uart_tx_en      <= 1'b0;
        uart_fft_over   <= 1'b0;
        rd_en           <= 1'b0;
        header_data_reg <= 8'h00;
    end else begin
        // Ĭ�Ͻ������ź�����
        rd_en      <= 1'b0;
        uart_tx_en <= 1'b0;

        // FSM ״̬ת��
        case (state_reg)
            // 0: ����״̬
            S_IDLE: begin
                count_reg <= 11'd0; // �������ݼ�����
                
                // ���FIFO���Ƿ������ݣ����У���ʼ����
                if (!rd_empty) begin
                    uart_fft_over   <= 1'b0; // �����һ֡����ɱ�־
                    header_data_reg <= 8'h05; // Ԥ���ص�һ��֡ͷ
                    state_reg       <= S_SEND_HEADER1; 
                end else begin
                    // ���ֿ��У��ȴ�����
                    state_reg       <= S_IDLE;
                end
            end
            
            // 1: ����֡ͷ1 (0x05)
            S_SEND_HEADER1: begin
                uart_tx_en   <= 1'b1; // ����ʹ�� (��ʱ uart_tx_data = 8'h05)
                state_reg    <= S_WAIT_HEADER1;
            end
            
            // 2: �ȴ�֡ͷ1�������
            S_WAIT_HEADER1: begin
                if (uart_tx_done) begin
                    header_data_reg <= 8'h64; // Ԥ���صڶ���֡ͷ
                    state_reg       <= S_SEND_HEADER2; 
                end else begin
                    state_reg       <= S_WAIT_HEADER1; // �����ȴ�
                end
            end

            // 3: ����֡ͷ2 (0x64)
            S_SEND_HEADER2: begin
                uart_tx_en   <= 1'b1; // ����ʹ�� (��ʱ uart_tx_data = 8'h64)
                state_reg    <= S_WAIT_HEADER2;
            end
            
            // 4: �ȴ�֡ͷ2�������
            S_WAIT_HEADER2: begin
                if (uart_tx_done) begin
                    // ֡ͷ������ϣ�׼����ʼ��������
                    // �ٴμ��FIFOȷ����ȫ
                    if (!rd_empty) begin
                        state_reg <= S_READ_FIFO;
                    end else begin
                        state_reg <= S_IDLE; // �쳣��FIFO���ˣ�����IDLE
                    end
                end else begin
                    state_reg <= S_WAIT_HEADER2; // �����ȴ�
                end
            end
            
            // 5: ��FIFO��ȡ����
            S_READ_FIFO: begin
                rd_en     <= 1'b1; // ����һ��ʱ�����ڵĶ�ʹ��
                state_reg <= S_SEND_UART; // ��һ��ȥ����
            end

            // 6: ����FIFO����
            S_SEND_UART: begin
                // (��ʱ uart_tx_data = rd_data, �� assign ��䴦��)
                uart_tx_en   <= 1'b1; // ����ʹ��
                state_reg    <= S_WAIT_UART;
            end

            // 7: �ȴ�UART���ݷ������
            S_WAIT_UART: begin
                if (uart_tx_done) begin
                    // ����Ƿ������һ������
                    if (count_reg == 11'd2047) begin // (0 �� 2047 �� 2048��)
                        state_reg <= S_FINISH;
                    end else begin
                        // ��δ���꣬׼������һ��
                        count_reg <= count_reg + 1;
                        if (!rd_empty) begin
                            state_reg <= S_READ_FIFO; // ��ȥ����һ������
                        end else begin
                            // ���󣺷���FIFOǷ�� (Underrun)
                            state_reg <= S_IDLE; 
                        end
                    end
                end else begin
                    // ���ڻ�û���꣬�����ȴ�
                    state_reg <= S_WAIT_UART;
                end
            end

            // 8: ���
            S_FINISH: begin
                uart_fft_over <= 1'b1; // ��λ��ɱ�־
                state_reg     <= S_IDLE; // �ص�IDLE״̬���ȴ���һ֡
            end

            default: begin
                state_reg <= S_IDLE;
            end
        endcase
    end
end

endmodule