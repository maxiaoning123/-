//���ֵ����ģ��
module vpp_measure(   
    input               rst_n,      // ��λ�ź�
    
    input               ad_clk,     // ADʱ��
    input      [7:0]    ad_data,    // AD��������
    input               ad_pulse,   // ��AD���εõ��������ź�
    output reg [7:0]    ad_vpp,     // AD���ֵ
    output reg [7:0]    ad_max,     // AD���ֵ
    output reg [7:0]    ad_min      // AD��Сֵ
);

//reg define
reg         vpp_flag;               // �������ֵ��־�ź�
reg         vpp_flag_d;             // vpp_flag ��ʱ
reg [7:0]   ad_data_max;            // ADһ�������ڵ����ֵ
reg [7:0]   ad_data_min;            // ADһ�������ڵ���Сֵ

//wire define
wire        vpp_flag_pos;           // vpp_flag�����ر�־�ź�
wire        vpp_flag_neg;           // vpp_flag�½��ر�־�ź�

//���ؼ�⣬�����ź�����/�½���
assign vpp_flag_pos = (~vpp_flag_d) & vpp_flag;
assign vpp_flag_neg = vpp_flag_d & (~vpp_flag);

//����vpp_flag��־һ������ʱ������
always @(posedge ad_pulse or negedge rst_n) begin
    if(!rst_n)
        vpp_flag <= 1'b0; 
    else 
        vpp_flag <= ~vpp_flag; 
end

//��vpp_flag��ʱһ��ADʱ������
always @(posedge ad_clk or negedge rst_n) begin
    if(!rst_n)
        vpp_flag_d <= 1'b0; 
    else 
        vpp_flag_d <= vpp_flag; 
end

//ɸѡһ������ʱ�������ڵ����/��Сֵ
always @(posedge ad_clk or negedge rst_n) begin
    if(!rst_n) begin
        ad_data_max <= 8'd0; 
        ad_data_min <= 8'd0;
    end
    else if(vpp_flag_pos)begin      //����ʱ�����ڿ�ʼʱ�Ĵ�AD����
        ad_data_max <= ad_data; 
        ad_data_min <= ad_data;
    end
    else if(vpp_flag_d) begin   
        if(ad_data > ad_data_max)
            ad_data_max <= ad_data; //�������ֵ
        if(ad_data < ad_data_min)
            ad_data_min <= ad_data; //������Сֵ
    end    
end

//���㱻��ʱ�������ڵķ��ֵ
always @(posedge ad_clk or negedge rst_n) begin
    if(!rst_n) begin
        ad_vpp <= 8'd0;
        ad_max <= 8'd0;
        ad_min <= 8'd0;
    end
    else if(vpp_flag_neg) begin
        ad_vpp <= ad_data_max - ad_data_min;
        ad_max <= ad_data_max;
        ad_min <= ad_data_min;
    end
end

endmodule