module auto_check(
    input         clk,
    input         rst_n,
    input         Goal_inc,//Ŀ��Ƶ�����Ӱ���
    input         Goal_dec,//Ŀ��Ƶ�ʼ�С����
    input [19:0]  ad_freq, // ʵ�ʲ�����Ƶ�ʣ���λ��Hz��
    
    output        Goal_flag // Ŀ��Ƶ���Ƿ��ڷ�Χ��
   );

// ------------------------------------------
// I. �������� (����Ƶ�ʵ�λ�� Hz)
// ------------------------------------------
localparam FREQ_RANGE_HZ    = 20'd1000;    // max��min֮��Ĺ̶���ֵ��1000 Hz
localparam ADJUST_STEP_HZ   = 20'd10000;   // ÿ������/���ٵĲ���ֵ��10 kHz (10000 Hz)

// Ƶ�����ƣ��������Ƶ�ʲ����� 1MHz, �� 1,000,000 Hz��
localparam MAX_LIMIT_HZ     = 20'd1000000; // 1MHz
localparam MIN_LIMIT_HZ     = 20'd10000;   // 10kHz

// ------------------------------------------
// II. �ڲ��źźͼĴ���
// ------------------------------------------
reg [19:0]    Goal_freq_max; // Ŀ��Ƶ�ʷ�Χ����
reg [19:0]    Goal_freq_min; // Ŀ��Ƶ�ʷ�Χ����

// ����ͬ���ͱ��ؼ�⣨�򻯴���ʵ���н���ʹ�ø����Ƶ������߼���
reg           Goal_inc_d;
reg           Goal_dec_d;
wire          inc_pulse;
wire          dec_pulse;

// ------------------------------------------
// III. ������������ (��Ϊ�����ؼ��)
// ------------------------------------------
always @(posedge clk or negedge rst_n) begin
    if (rst_n == 1'b0) begin
        Goal_inc_d <= 1'b0;
        Goal_dec_d <= 1'b0;
    end else begin
        Goal_inc_d <= Goal_inc;
        Goal_dec_d <= Goal_dec;
    end
end

assign inc_pulse = Goal_inc & (~Goal_inc_d); // ���Ӱ�����������
assign dec_pulse = Goal_dec & (~Goal_dec_d); // ��С������������

// ------------------------------------------
// IV. Ŀ��Ƶ�ʼĴ��������߼�
// ------------------------------------------
always @(posedge clk or negedge rst_n) begin
    if (rst_n == 1'b0) begin
        // ��λʱ��ʼ��Ŀ��Ƶ�ʷ�Χ (����� 10kHz ��ʼ)
        Goal_freq_min <= 20'd10000; 
        Goal_freq_max <= 20'd10000 + FREQ_RANGE_HZ; // 11kHz
    end else if (inc_pulse) begin
        // Ŀ��Ƶ������
        // ��� Goal_freq_max ���Ӻ��Ƿ񳬹��������
        if (Goal_freq_max + ADJUST_STEP_HZ <= MAX_LIMIT_HZ) begin
            Goal_freq_min <= Goal_freq_min + ADJUST_STEP_HZ;
            Goal_freq_max <= Goal_freq_max + ADJUST_STEP_HZ;
        end else begin
            // �ﵽ���ޣ����ֲ���
            Goal_freq_min <= Goal_freq_min; 
            Goal_freq_max <= Goal_freq_max;
        end
    end else if (dec_pulse) begin
        // Ŀ��Ƶ�ʼ�С
        // ��� Goal_freq_min ��С���Ƿ������С����
        if (Goal_freq_min >= MIN_LIMIT_HZ + ADJUST_STEP_HZ) begin 
            Goal_freq_min <= Goal_freq_min - ADJUST_STEP_HZ;
            Goal_freq_max <= Goal_freq_max - ADJUST_STEP_HZ;
        end else begin
            // �ﵽ���ޣ����ֲ���
            Goal_freq_min <= Goal_freq_min; 
            Goal_freq_max <= Goal_freq_max;
        end
    end
    // ע�⣺���� Goal_freq_max �� Goal_freq_min ����ͨ���Ӽ� ADJUST_STEP_HZ ������
    // �ҳ�ʼֵ���� Goal_freq_max = Goal_freq_min + FREQ_RANGE_HZ��
    // ����֮��Ĳ�ֵ (FREQ_RANGE_HZ) ���Զ����ֲ��䡣
end

// ------------------------------------------
// V. Ŀ��Ƶ�ʼ���߼�
// ------------------------------------------
assign Goal_flag = (ad_freq >= Goal_freq_min) && (ad_freq <= Goal_freq_max);

endmodule