/*
 * ģ����: wave_detector_auto (�Կز�����)
 * ��  ��: ��Ⲩ�������Ҳ����Ƿ����������п��Ʋ������ڡ�
 * ʱ  ��: ad_clk �������ݲ������߼�ִ�С�
 */
module wave_detector (
    input             clk,         // AD����ʱ�ӣ���ad_clk
    input             rst_n,       // ϵͳ��λ
    input      [7:0]  ad_data_in,  // �����ƽ����AD���� (ad_avg_data)
    input      [7:0]  ad_max_in,   // 8λ��ĵ�ǰ�������ֵ
    input      [7:0]  ad_min_in,   // 8λ��ĵ�ǰ������Сֵ
    output reg        is_square    // ʶ������1'b1 = ������1'b0 = ���Ҳ�
);

// --- �������� ---
// �����жϵ���ֵ
parameter THRESHOLD_CNT = 10; 

// �ڲ���̬��ֵ����
// UPPER_THRESH_DYN = ad_max_in - 10
// LOWER_THRESH_DYN = ad_min_in + 10

// --- ״̬������ ---
localparam S_WAIT_LOW  = 2'd0; // �ȴ����ݵ��� LOWER_THRESH_DYN
localparam S_COUNT_UP  = 2'd1; // ������������ֵ֮��仯ʱ����
localparam S_WAIT_HIGH = 2'd2; // �ȴ����ݸ��� UPPER_THRESH_DYN

// --- �ڲ��ź� ---
reg  [15:0] count/* synthesis PAP_MARK_DEBUG="1"*/;         // �����������ڼ�¼��������ʱ������
reg  [1:0]  state/* synthesis PAP_MARK_DEBUG="1"*/;         // ״̬���Ĵ���

// ���㶯̬��ֵ
// ȷ�������ͼӷ���������������� 8 λ���Ͽ����Խ�С
wire [7:0] UPPER_THRESH_DYN;
wire [7:0] LOWER_THRESH_DYN;

// ��̬������ֵ��ad_max_in - 10 �� ad_min_in + 10
// ʹ�����������ȷ����ֵ�������磬ad_max_in - 10 ����Ϊ 10��
assign UPPER_THRESH_DYN = (ad_max_in > 8'd10) ? (ad_max_in - 8'd10) : 8'd10; 
assign LOWER_THRESH_DYN = (ad_min_in < 8'd245) ? (ad_min_in + 8'd10) : 8'd245;

// --- ��������״̬���߼� ---
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        state     <= S_WAIT_LOW;
        count     <= 16'd0;
        is_square <= 1'b0; // Ĭ�����Ҳ�
    end else begin
        case (state)
            S_WAIT_LOW: begin
                // ״̬0���ȴ������½��� LOWER_THRESH_DYN ����
                if (ad_data_in < LOWER_THRESH_DYN) begin
                    // �Ѿ�������ֵ��׼����ʼ�����ؼ���
                    state <= S_COUNT_UP;
                    count <= 16'd0; // ���ü�����
                end
            end
            
            S_COUNT_UP: begin
                // ״̬1����ʼ������ֱ�����δﵽ UPPER_THRESH_DYN
                if (ad_data_in < LOWER_THRESH_DYN) begin
                    // ������������½������»ص��ȴ���λ״̬�����ü���
                    state <= S_WAIT_LOW;
                    count <= 16'd0;
                end else if (ad_data_in >= UPPER_THRESH_DYN) begin
                    // �ﵽ��ֵ�����������
                    state <= S_WAIT_HIGH;
                    
                    // --- �о��߼� ---
                    if (count <= THRESHOLD_CNT) begin
                        // ������С������ǳ��� -> ����
                        is_square <= 1'b1;
                    end else begin
                        // �����ϴ󣬱仯ƽ�� -> ���Ҳ�
                        is_square <= 1'b0;
                    end
                end else begin
                    // �������������У���������
                    count <= count + 1'b1;
                    // ������������
                    if (count == 16'hFFFF) begin 
                         state <= S_WAIT_HIGH; 
                         is_square <= 1'b0; // �仯̫������Ϊ���Ҳ�
                    end
                end
            end
            
            S_WAIT_HIGH: begin
                // ״̬2���ȴ������½��� LOWER_THRESH_DYN ���£��Կ�ʼ��һ���ж�
                if (ad_data_in < LOWER_THRESH_DYN) begin
                    state <= S_WAIT_LOW;
                end
            end
            
            default: state <= S_WAIT_LOW;
        endcase
    end
end

endmodule