module avg_filter_8bit #(
    parameter N = 16  // ƽ��������2���ݴΣ���2/4/8/16��NԽ���˲�Խǿ��
) (
    input               clk,        // ������AD����ʱ�ӣ���ad_clk��
    input               rst_n,      // �͵�ƽ��Ч��λ
    input  [7:0]        data_in,    // 8bit ADԭʼ����
    output reg [7:0]    data_out    // 8bit �˲�������
);

// �ۼӺ�λ��8bit + log2(N)�������������N=8ʱ��11bit��
reg [7 + $clog2(N):0] sum;
reg [7:0] buf1 [N-1:0];  // �������ڻ���
integer i;

always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        sum <= 0;
        data_out <= 0;
        for (i = 0; i < N; i = i + 1) buf1[i] <= 0;
    end else begin
        // �Ƴ�������ݣ����������
        sum <= sum - buf1[N-1] + data_in;
        // ������λ
        for (i = N-1; i > 0; i = i - 1) buf1[i] <= buf1[i-1];
        buf1[0] <= data_in;
        // ��λ���������NΪ2���ݴΣ�Ч����ߣ�
        data_out <= sum >> $clog2(N);
    end
end

endmodule