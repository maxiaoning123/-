module median_filter_8bit #(
    parameter WINDOW = 3  // ���ڴ�С��3/5/7��������3����ʡ��Դ��
) (
    input               clk,
    input               rst_n,
    input  [7:0]        data_in,
    output reg [7:0]    data_out
);

reg [7:0] buf1 [WINDOW-1:0];  // �������ڻ���
reg [7:0] temp [WINDOW-1:0]; // ������ʱ����
integer i, j;

always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        for (i = 0; i < WINDOW; i = i + 1) buf1[i] <= 0;
        data_out <= 0;
    end else begin
        // ������λ���Ƴ�������ݣ�����������
        for (i = WINDOW-1; i > 0; i = i - 1) buf1[i] <= buf1[i-1];
        buf1[0] <= data_in;
        
        // �������ݵ���ʱ���飨�����޸�ԭ���棩
        for (i = 0; i < WINDOW; i = i + 1) temp[i] <= buf1[i];
        
        // ð������8bit��������Ч�ʸߣ�
        for (i = 0; i < WINDOW-1; i = i + 1) begin
            for (j = 0; j < WINDOW-1 - i; j = j + 1) begin
                if (temp[j] > temp[j+1]) begin
                    temp[j] <= temp[j+1];
                    temp[j+1] <= temp[j];
                end
            end
        end
        
        // ȡ�м�ֵ������Ϊ������ֱ��ȡ�м�������
        data_out <= temp[WINDOW/2];
    end
end

endmodule