module measure(
    input               clk_50M ,       // ʱ��
    input               rst_n  ,    // ��λ�ź�

    input                ad_clk,     // ADʱ��
    input      [7:0]     ad_data_in,
    output [31:0]        duty,
    output [19:0]        ad_freq,
    output [7:0]         ad_max,
    output [7:0]         ad_min
    

    
);
wire              ad_pulse/* synthesis PAP_MARK_DEBUG="1"*/;   //pulse_genģ������������ź�,�����ڵ���
wire              ad_pulse_reg/* synthesis PAP_MARK_DEBUG="1"*/;   

wire  [7:0]    ad_vpp;   // AD���ֵ 

//wire      [7:0]    ad_min;      // AD��Сֵ
//parameter define
parameter CLK_FS = 26'd50_000_000;  // ��׼ʱ��Ƶ��ֵ

//wire clk_100m;
wire [17:0]o_duty_num;

signal_fir u_signal_fir(
    .sys_clk       (clk_50M),     // ����ϵͳʱ�ӣ�ȷ���˲�ʱ����ϵͳͬ����
    .rst_n         (rst_n),   // ����ϵͳ��λ���͵�ƽ��Ч��
    .TTL_signal    (ad_pulse_reg),     // �����ë�̵�ԭʼTTL�ź�
    .TTL_signal_fir(ad_pulse) // ����˲�����ȶ�TTL�ź�
);


//��������ģ��
pulse_gen u_pulse_gen(
    .rst_n          (rst_n),        //ϵͳ��λ���͵�ƽ��Ч

    .trig_level     (8'd128),   // ������ƽ
    .ad_clk         (ad_clk),       //AD9280����ʱ��
    .ad_data        (ad_data_in),      //AD��������

    .ad_pulse       (ad_pulse_reg)      //����������ź�
    );

//�Ⱦ���Ƶ�ʼ�ģ��
cymometer #(
    .CLK_FS         (CLK_FS)        // ��׼ʱ��Ƶ��ֵ
) u_cymometer(
    .clk_fs         (clk_50M),
    .rst_n          (rst_n),

    .clk_fx         (ad_pulse),     // ����ʱ���ź�
    .data_fx        (ad_freq)       // ����ʱ��Ƶ�����
    );

//������ֵ
vpp_measure u_vpp_measure(
    .rst_n          (rst_n),
    
    .ad_clk         (ad_clk), 
    .ad_data        (ad_data_in),
    .ad_pulse       (ad_pulse),
    .ad_vpp         (ad_vpp),
    .ad_max         (ad_max),
    .ad_min         (ad_min)
    );
wire [31:0]high_time;
wire [31:0]low_time;

duty_cycle u_duty_cycle(
    .clk(clk_50M),
    
    .rst_n(rst_n),
    .signal_in(ad_pulse),
    .high_time(high_time),
    .low_time(low_time),
    .duty(duty)
);
endmodule
