module top(
    input                     clk_27M,//27m Hz
    input                     rst,
    input                     key_add_1000hz,
    input                     key_add_10hz,
    input                     key_inc_duty,         // ռ�ձ����Ӱ���
    input                     key_dec_duty,         // ռ�ձȼ��ٰ���
    input                     key_change_wave,      // �����л�����
    input            		  uart_rxd /* synthesis PAP_MARK_DEBUG="1"*/,   
    output           		  uart_txd /* synthesis PAP_MARK_DEBUG="1"*/,
    input            		  uart_rxd1 /* synthesis PAP_MARK_DEBUG="1"*/,   
    output           		  uart_txd1 /* synthesis PAP_MARK_DEBUG="1"*/,
    output        wire        da_clk /* synthesis PAP_MARK_DEBUG="1"*/,
    output        wire        ad_clk /* synthesis PAP_MARK_DEBUG="1"*/,
    output        wire [7:0]  da_data /* synthesis PAP_MARK_DEBUG="1"*/,
    input         wire [7:0]  ad_data_in/* synthesis PAP_MARK_DEBUG="1"*/,
    
    output        wire        auto_check_led,
    output        wire        led_wave,
    output                    lcd_spi_sclk    ,// ��Ļspiʱ�ӽӿ�
    output                    lcd_spi_mosi    ,// ��Ļspi���ݽӿ�
    output                    lcd_spi_cs      ,// ��Ļspiʹ�ܽӿ�     
    output                    lcd_dc          ,// ��Ļ ����/���� �ӿ�
    output                    lcd_reset       ,// ��Ļ��λ�ӿ�
    output                    lcd_blk          // ��Ļ����ӿ� 
   );

//key signals
wire key_add_1000hz_neg;  // Ƶ��+1000Hz�����������½���
wire key_add_10hz_neg;    // Ƶ��+10Hz�����������½���
wire key_inc_duty_neg;    // ռ�ձ����Ӱ����������½���
wire key_dec_duty_neg;    // ռ�ձȼ��ٰ����������½���
wire key_change_wave_neg; // �����л������������½���

//DDS signals
wire [7:0]    square_out/* synthesis PAP_MARK_DEBUG="1"*/; //��������
wire [7:0]    sin_out/* synthesis PAP_MARK_DEBUG="1"*/;    //���Ҳ�����
wire          wave_flag/* synthesis PAP_MARK_DEBUG="1"*/;  //���������־ 0�����Ҳ� 1������ Ĭ��Ϊ0
//measure signals
wire [31:0]        duty       ;
wire [19:0]        ad_freq    ;
wire [7:0]         ad_max     ;
wire [7:0]         ad_min     ;
//fir signals
wire  [7:0]  ad_avg_data/* synthesis PAP_MARK_DEBUG="1"*/;
//fft signals
wire         fft_over/* synthesis PAP_MARK_DEBUG="1"*/;
wire         fft_start/* synthesis PAP_MARK_DEBUG="1"*/;
wire         lcd_draw_over/* synthesis PAP_MARK_DEBUG="1"*/;
wire [7:0]   o_fft_data_re/* synthesis PAP_MARK_DEBUG="1"*/;
wire [7:0]   o_fft_data_im/* synthesis PAP_MARK_DEBUG="1"*/;
wire         o_fft_data_vaild/* synthesis PAP_MARK_DEBUG="1"*/;
wire [31:0]  o_fft_data;
wire [7:0]   fft_data/* synthesis PAP_MARK_DEBUG="1"*/;

//pll signals
wire pll_lock;
wire pll1_lock;
wire clk_50M;
wire clk_30M;
wire rst_n;
//uart
wire            uart_tx_en; 
wire            uart_rx_done; 
wire            uart_tx_done; 
wire  [7:0]     uart_tx_data; 
wire  [7:0]     uart_rx_data; 
wire            uart_fft_over;
//auto check signals
wire         Goal_inc/* synthesis PAP_MARK_DEBUG="1"*/;
wire         Goal_dec/* synthesis PAP_MARK_DEBUG="1"*/;
assign rst_n = rst && pll_lock && pll1_lock ;
assign da_clk = ~ad_clk;
assign da_data = wave_flag ? square_out : sin_out;

pll_30m u_pll1 (
  .clkout0(clk_30M),    // output
  .lock(pll1_lock),          // output
  .clkin1(clk_27M)       // input
);
pll u_pll (
  .clkout0(ad_clk),    // output
  .clkout1(clk_50M),    // output
  .lock(pll_lock),          // output
  .clkin1(clk_30M)       // input
);


DDS_wave u_DDS_wave(
    .clk            (clk_50M),         // ����DDS����ʱ��
    .rst_n          (rst_n),       // ����ϵͳ��λ
    .key_add_1000hz (key_add_1000hz_neg),  // �����������+1000Hz����
    .key_add_10hz   (key_add_10hz_neg),    // �����������+10Hz����
    .key_inc_duty   (key_inc_duty_neg),    // �����������ռ�ձ����Ӱ���
    .key_dec_duty   (key_dec_duty_neg),    // �����������ռ�ձȼ��ٰ���
    .key_change_wave(key_change_wave_neg), // ����������Ĳ����л�����
    .wave_flag      (wave_flag),       //���������־ 0�����Ҳ� 1������ Ĭ��Ϊ0 
    .square_data    (square_out),      // �������
    .sin_data       (sin_out)          // ���Ҳ����
);


measure u_measure (
    // ����˿�����
    .clk_50M      (clk_50M),    // ����ϵͳ50MHzʱ��
    .rst_n        (rst_n),      // ����ϵͳ��λ�ź�
    .ad_data_in   (ad_avg_data),     // �����ⲿAD��������
    .ad_clk       (ad_clk),         // ���ADʱ�ӣ���ֱ�����ӵ�ADоƬ��ʱ�����ţ�
    // ����˿�����
    
    .duty         (duty),     // ռ�ձȽ�����
    .ad_freq      (ad_freq),        // Ƶ�ʽ�����
    .ad_max       (ad_max),          // ���ֵ������
    .ad_min       (ad_min)
);

auto_check u_auto_check (
    .clk        ( clk_50M          ), // ���룺ϵͳʱ��
    .rst_n      ( rst_n        ), // ���룺��λ�ź� (����Ч)
    .Goal_inc   ( Goal_inc        ), // ���룺Ŀ��Ƶ�����Ӱ���
    .Goal_dec   ( Goal_dec        ), // ���룺Ŀ��Ƶ�ʼ�С����
    .ad_freq    ( ad_freq    ), // ���룺ʵ�ʲ�����Ƶ��ֵ [19:0]
    
    .Goal_flag  ( auto_check_led    )  // �����ʵ��Ƶ���Ƿ���Ŀ�귶Χ��
);

wave_detector u_wave_detector (
    .clk          (ad_clk),         // ����AD����ʱ��
    .rst_n        (rst_n),
    .ad_data_in   (ad_avg_data),    // ����ƽ�����AD����
    .ad_max_in    (ad_max),         // ���Ӳ���ģ������� Max
    .ad_min_in    (ad_min),         // ���Ӳ���ģ������� Min
    .is_square    (led_wave)
);

bluetooth_data u_bluetooth_data (
    .clk            (clk_50M),
    .ad_clk         (ad_clk),
    .rst_n          (rst_n),
    .fft_data       (fft_data),
    .fft_data_vaild (o_fft_data_vaild),
    .uart_tx_done   (uart_tx_done),
    .uart_tx_en     (uart_tx_en),
    .uart_tx_data   (uart_tx_data),
    .uart_fft_over  (uart_fft_over)
);

uart_top uart2_top_inst (
    .sys_clk      (clk_50M),    // ϵͳʱ�ӣ����� UART �ڲ�����������
    .sys_rst_n    (rst_n),        // ϵͳ��λ���͵�ƽ��Ч����ģ�鶨��һ�£�
    
    .uart_rxd     (uart_rxd1), // �����ⲿ UART ��������
    .uart_txd     (uart_txd1), // �����ⲿ UART ��������
    
    .uart_tx_en   (uart_tx_en),   
    .uart_rx_done (uart_rx_done), 
    .uart_tx_done (uart_tx_done), 
    
    .uart_tx_data (uart_tx_data), 
    .uart_rx_data (uart_rx_data)  
);



fft_lcd_state_control u_fft_lcd_state_control(
    .clk        (ad_clk),     
    .rst_n      (rst_n),   // ��λ�źţ�����Ч��
    .lcd_draw_over(uart_fft_over),
    .ad_data    (ad_avg_data),     // AD�ɼ���������
    .fft_over   (fft_over),    // FFT��������ź�����
    .fft_start  (fft_start)    // FFT�����ź����
);


fft_control u_fft_control (
    .clk            (ad_clk),      
    .rst_n          (rst_n),    // ����ϵͳ��λ
    .fft_start      (fft_start),
    .fft_over       (fft_over),
    .i_fft_data     (ad_avg_data),      // ������������
    .fft_data       (fft_data),
    .o_fft_data     (o_fft_data),
    .o_fft_data_vaild(o_fft_data_vaild),
    .o_fft_data_re     (o_fft_data_re),  // �����������
    .o_fft_data_im     (o_fft_data_im)
);

lcd_top u_lcd_top(
    .sys_clk         (clk_50M   ),  // ����ϵͳʱ��
    .sys_rst_n       (rst_n     ),  // ����ϵͳ��λ
    .ad_clk          (ad_clk   ), 
    .o_fft_data_vaild(o_fft_data_vaild), 
    .o_fft_data      (fft_data      ),
    .lcd_draw_over   (lcd_draw_over),
    // LCD��Ļ�ӿ�����
    .lcd_spi_sclk    (lcd_spi_sclk  ),
    .lcd_spi_mosi    (lcd_spi_mosi  ),
    .lcd_spi_cs      (lcd_spi_cs    ),
    .lcd_dc          (lcd_dc        ),
    .lcd_reset       (lcd_reset     ),
    .lcd_blk         (lcd_blk       )
);

Bluetooth_send u_Bluetooth_send(
    .sys_clk       (clk_50M),      // ����ϵͳʱ��
    .rst_n         (rst_n),    // ����ϵͳ��λ���͵�ƽ��Ч��
    
    .uart_rxd      (uart_rxd),// ��������ģ���UART���նˣ�FPGA�����������ݣ�
    .uart_txd      (uart_txd),// ��������ģ���UART���Ͷˣ�FPGA�������������ݣ�
    .Goal_inc      (Goal_inc), 
    .Goal_dec      (Goal_dec), 
    .duty_cycle    (duty),   // ����ռ�ձȲ�������
    .ad_fred       (ad_freq),      // ����Ƶ�ʲ������ݣ�����ԭ"ad_fred"ƴд��
    .ad_max        (ad_max)        // �������ֵ��������
);


avg_filter_8bit #(
    .N(16)  // �ɵ���Ϊ4/16��������������Ż�
) u_avg_filter (
    .clk(ad_clk),         // ����AD����ʱ�ӣ���ad_clk��
    .rst_n(rst_n), // ����ϵͳ��λ
    .data_in(ad_data_in), // ����8bit ADԭʼ����
    .data_out(ad_avg_data) // ���ƽ���������
);



key_debounce u_key_1000hz_debounce (
    .sys_clk       (clk_50M),         // ϵͳʱ������
    .rst_n         (rst_n),           // ��λ�źţ�����Ч��
    .key           (key_add_1000hz),  // ԭʼ�������루+1000Hz��
    .button_negedge(key_add_1000hz_neg) // ��������½����ź�
);

key_debounce u_key_10hz_debounce (
    .sys_clk       (clk_50M),         // ϵͳʱ������
    .rst_n         (rst_n),           // ��λ�źţ�����Ч��
    .key           (key_add_10hz),    // ԭʼ�������루+10Hz��
    .button_negedge(key_add_10hz_neg) // ��������½����ź�
);

key_debounce u_key_inc_duty_debounce (
    .sys_clk       (clk_50M),         // ϵͳʱ������
    .rst_n         (rst_n),           // ��λ�źţ�����Ч��
    .key           (key_inc_duty),    // ԭʼ�������루ռ�ձ�+��
    .button_negedge(key_inc_duty_neg) // ��������½����ź�
);


key_debounce u_key_dec_duty_debounce (
    .sys_clk       (clk_50M),         // ϵͳʱ������
    .rst_n         (rst_n),           // ��λ�źţ�����Ч��
    .key           (key_dec_duty),    // ԭʼ�������루ռ�ձ�-��
    .button_negedge(key_dec_duty_neg) // ��������½����ź�
);



key_debounce u_key_change_wave_debounce (
    .sys_clk       (clk_50M),         // ϵͳʱ������
    .rst_n         (rst_n),           // ��λ�źţ�����Ч��
    .key           (key_change_wave),     // ԭʼ�������루�л���
    .button_negedge(key_change_wave_neg)  // ��������½����ź�
);




endmodule
