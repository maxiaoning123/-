module pulse_gen(
    input           rst_n,      //ϵͳ��λ���͵�ƽ��Ч
    
    input  [7:0]    trig_level,
    input           ad_clk,     //AD����ʱ��
    input  [7:0]    ad_data,    //AD��������
    
    output          ad_pulse    //����������ź�
);

parameter THR_DATA = 3;

//reg define
reg          pulse;
reg          pulse_delay;

assign ad_pulse = pulse & pulse_delay;

//���ݴ�����ƽ���������AD����ֵת���ɸߵ͵�ƽ
always @ (posedge ad_clk or negedge rst_n)begin
    if(!rst_n)
        pulse <= 1'b0;
    else begin
        if((trig_level >= THR_DATA) && (ad_data < trig_level - THR_DATA))
            pulse <= 1'b0;
        else if(ad_data > trig_level + THR_DATA)
            pulse <= 1'b1;
    end    
end

//��ʱһ��ʱ�����ڣ�������������
always @ (posedge ad_clk or negedge rst_n)begin
    if(!rst_n)
        pulse_delay <= 1'b0;
    else
        pulse_delay <= pulse;
end

endmodule