module kalman_filter_8bit (
    input               clk,
    input               rst_n,
    input  [7:0]        data_in,    // 8bit AD����
    output reg [7:0]    data_out    // 8bit �˲����
);

// 8bit���������Q=����������R=�۲���������΢����
parameter Q = 8'd2;    // ����������ԽСԽ������ʷֵ���˲�Խƽ����
parameter R = 8'd10;   // �۲�������ԽСԽ����AD���ݣ���ӦԽ�죩

reg [15:0] P = 16'd0;  // Э�����չλ����������
reg [15:0] LastP = 16'd0;
reg [15:0] Kg = 16'd0; // ���������棨16λ����������8λ����+��8λС����
reg [7:0] LastOut = 8'd0;

always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        P <= 16'd0;
        LastP <= 16'd0;
        Kg <= 16'd0;
        LastOut <= 8'd0;
        data_out <= 8'd0;
    end else begin
        // Ԥ��Э����
        P <= LastP + Q;
        // ���㿨�������棨���������㣬���⸡������
        Kg <= (P << 8) / (P + R);  // ����8λ�Ŵ�����8λ��ԭ
        // ���Ź��ƣ����������
        if (data_in > LastOut) begin
            data_out <= LastOut + ((Kg * (data_in - LastOut)) >> 8);
        end else begin
            data_out <= LastOut - ((Kg * (LastOut - data_in)) >> 8);
        end
        // ����Э����
        LastP <= ((16'd255 - Kg[15:8]) * P) >> 8;  // ȡKg��������
        LastOut <= data_out;
    end
end

endmodule